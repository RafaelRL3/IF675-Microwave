module encoder (
    input wire [8:0]keypad,
    input wire clock,
    input wire enable, 
    output wire [3:0]D,
    output wire pgt_1Hz,
    output wire loadn
);

    
endmodule